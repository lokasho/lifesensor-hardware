.title KiCad schematic
R3 "/ecginputprotection/in2_LA" "/in_LA" 10k
R7 "/ecginputprotection/neon_LA" /ecginputprotection/in2_LA" 10k
V1 /in_LA GNDPWR pulse(0 4.8k 0 10u 10m 10u)
.tran 10u 20m 0 
.end
